//------------------------------------------------
// Nguyen Van Chuyen
// 2023-12-14
//
//
//-------------------------------------------------
//
// Class Description
//
////////////////////////////////////////////////////

package env_pkg;

  // Standard UVM import & include:
import uvm_pkg::*;
`include "uvm_macros.svh"

import add_agent_pkg::*;
import mul_agent_pkg::*;


  // Includes:
  `include "vsequencer.svh"
  `include "sco.svh"
  `include "env.svh"

endpackage: env_pkg
