//------------------------------------------------
// Nguyen Van Chuyen
// 2023-12-22s
//
//
//-------------------------------------------------
//
// Class Description


`ifndef MUL_AGENT_PKG_SV
`define MUL_AGENT_PKG_SV

package mul_agent_pkg;
	
import uvm_pkg::*;
`include "uvm_macros.svh"

`include "mul_transaction.svh"
`include "mul_driver.svh"
`include "mul_mon.svh"
`include "mul_agent.svh"


endpackage : mul_agent_pkg

`endif

