//------------------------------------------------
// Nguyen Van Chuyen
// 2023-12-22s
//
//
//-------------------------------------------------
//
// Class Description


`ifndef ADD_AGENT_PKG_SV
`define ADD_AGENT_PKG_SV

package add_agent_pkg;
	
import uvm_pkg::*;
`include "uvm_macros.svh"

`include "add_transaction.svh"
`include "add_driver.svh"
`include "add_mon.svh"
`include "add_agent.svh"

endpackage : add_agent_pkg

`endif

